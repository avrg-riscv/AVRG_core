//this is a interface example
